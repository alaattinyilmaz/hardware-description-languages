// `timescale 1ns / 1ps
module intra_predictor (I, J, K, L, M, N, O, P, a1,a2,a3,a4,b1,b2,b3,b4,c1,c2,c3,c4,d1,d2,d3,d4);
input [7:0] I, J, K, L, M, N, O, P;
output reg [7:0] a1,a2,a3,a4,b1,b2,b3,b4,c1,c2,c3,c4,d1,d2,d3,d4;
reg [17: 0] temp;

always @ *
begin

//////////////////////

temp = ( ( (I << 4) + (I << 3) + (I << 2) + I ) + ( (J << 7) + (J << 6) + (J << 5) + (J << 3) + (J << 2) ) - ( (K << 3) + K ) ) >> 8;
a1 = temp;

temp = ( ( (J << 5) + (J << 4) + (J << 3) + (J << 2) + J ) - ( (I << 3) + I ) + ( (K << 7) + (K << 6) + (K << 4) + (K << 3) + K ) - ( (L << 3) + (L << 2) + L ) ) >> 8;
a2 = temp;

temp = ( ( (K << 6) + (K << 4) + (K << 3) + K ) - ( (J << 3) + (J << 2) ) + ( (L << 7) + (L << 6) + (L << 1) + L ) - (M << 4) ) >> 8;
a3 = temp;

temp = ( ( (L << 6) + (L << 5) + (L << 4) + (L << 2) ) - ( (K << 3) + (K << 2) + (K << 1) ) + ( (M << 7) + (M << 4) + (M << 3) + (M << 1) ) ) >> 8;
a4 = temp;


//////////////////////

temp = ( ( (J << 4) + (J << 3) + (J << 2) + J ) + ( (K << 7) + (K << 6) + (K << 5) + (K << 3) + (K << 2) ) - ( (L << 3) + L ) ) >> 8;
b1 = temp;

temp = ( ( (K << 5) + (K << 4) + (K << 3) + (K << 2) + K ) - ( (J << 3) + J ) + ( (L << 7) + (L << 6) + (L << 4) + (L << 3) + L ) - ( (M << 3) + (M << 2) + M ) ) >> 8;
b2 = temp;

temp = ( ( (L << 6) + (L << 4) + (L << 3) + L ) - ( (K << 3) + (K << 2) ) + ( (M << 7) + (M << 6) + (M << 1) + M ) - (N << 4) ) >> 8;
b3 = temp;

temp = ( ( (M << 6) + (M << 5) + (M << 4) + (M << 2) ) - ( (L << 3) + (L << 2) + (L << 1) ) + ( (N << 7) + (N << 4) + (N << 3) + (N << 1) ) ) >> 8;
b4 = temp;


//////////////////////

temp = ( ( (K << 4) + (K << 3) + (K << 2) + K ) + ( (L << 7) + (L << 6) + (L << 5) + (L << 3) + (L << 2) ) - ( (M << 3) + M ) ) >> 8;
c1 = temp;

temp = ( ( (L << 5) + (L << 4) + (L << 3) + (L << 2) + L ) - ( (K << 3) + K ) + ( (M << 7) + (M << 6) + (M << 4) + (M << 3) + M ) - ( (N << 3) + (N << 2) + N ) ) >> 8;
c2 = temp;

temp = ( ( (M << 6) + (M << 4) + (M << 3) + M ) - ( (L << 3) + (L << 2) ) + ( (N << 7) + (N << 6) + (N << 1) + N ) - (O << 4) ) >> 8;
c3 = temp;

temp = ( ( (N << 6) + (N << 5) + (N << 4) + (N << 2) ) - ( (M << 3) + (M << 2) + (M << 1) ) + ( (O << 7) + (O << 4) + (O << 3) + (O << 1) ) ) >> 8;
c4 = temp;


//////////////////////

temp = ( ( (L << 4) + (L << 3) + (L << 2) + L ) + ( (M << 7) + (M << 6) + (M << 5) + (M << 3) + (M << 2) ) - ( (N << 3) + N ) ) >> 8;
d1 = temp;

temp = ( ( (M << 5) + (M << 4) + (M << 3) + (M << 2) + M ) - ( (L << 3) + L ) + ( (N << 7) + (N << 6) + (N << 4) + (N << 3) + N ) - ( (O << 3) + (O << 2) + O ) ) >> 8;
d2 = temp;

temp = ( ( (N << 6) + (N << 4) + (N << 3) + N ) - ( (M << 3) + (M << 2) ) + ( (O << 7) + (O << 6) + (O << 1) + O ) - (P << 4) ) >> 8;
d3 = temp;

temp = ( ( (O << 6) + (O << 5) + (O << 4) + (O << 2) ) - ( (N << 3) + (N << 2) + (N << 1) ) + ( (P << 7) + (P << 4) + (P << 3) + (P << 1) ) ) >> 8;
d4 = temp;

end

endmodule